package shared_pkg ;

	logic test_finished ;
	integer error_count ;
	integer correct_count ;
	
endpackage 	